module adder (
    input  logic [3:0] a,
    input  logic [3:0] b,
    input  logic       carry_in,
    output logic [3:0] sum,
    output logic       carry_out
);


endmodule
