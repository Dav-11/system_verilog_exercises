`timescale 1ns / 10ps

module wb_mux_tb;

endmodule: wb_mux_tb
